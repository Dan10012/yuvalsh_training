




package enforcer_pack;
	
	typedef enum {
		WAIT_FOR_SOP,
		WAIT_FOR_EOP
	} enforcer_sm_t;



endpackage