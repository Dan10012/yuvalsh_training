if (
) begin
	/* code */
end